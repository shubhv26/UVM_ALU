
class scoreboard extends uvm_scoreboard;
  `uvm_component_utils(scoreboard)
  
  uvm_tlm_analysis_fifo#(seq_item)item_collected;
  seq_item seq;
  
    
  function new(string name,uvm_component parent);
    super.new(name,parent);
  endfunction:new
  
    //////////////////BUILD PHASE////////////////////
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    item_collected=new("items_collected",this);
  endfunction:build_phase
  
  
  ///////////// RUN PHASE////////////////////////////
  
  virtual task run_phase(uvm_phase phase);
    forever begin
      item_collected.get(seq);
      if(seq.sel== 3'b000)
        begin
        		if(seq.A+seq.B == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
          		`uvm_info(get_type_name(),$sformatf(" Value of SUM = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end
        
      else if(seq.sel==3'b001)
        begin
          if(seq.A+(~seq.B+1) == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
                `uvm_info(get_type_name(),$sformatf(" Value of DIFFERENCE = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end
        
      else if(seq.sel==3'b010)
        begin
          if(seq.A & seq.B == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
                `uvm_info(get_type_name(),$sformatf(" Value of A & B = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end
        
      else if(seq.sel==3'b011)
        begin
          		if(seq.A | seq.B == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
                `uvm_info(get_type_name(),$sformatf(" Value of A | B = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end
        
      else if(seq.sel== 3'b100)
        begin
          if(seq.A*seq.B == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
                `uvm_info(get_type_name(),$sformatf(" Value of PRODUCT = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end

      else if(seq.sel== 3'b101)
        begin
          if(seq.A ^ seq.B == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
            `uvm_info(get_type_name(),$sformatf(" Value of A xor B = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end
     
      else if(seq.sel== 3'b110)
        begin
          if(~(seq.A&seq.B) == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
            `uvm_info(get_type_name(),$sformatf(" Value of A nand B = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end
      
      else if(seq.sel== 3'b111)
        begin
          if(~(seq.A | seq.B) == seq.Result) begin
          	    $display("------------------------SCOREBOARD-----------------------------------------");
        		`uvm_info(get_type_name(),$sformatf(" TEST PASS "),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of A = %0d", seq.A),UVM_LOW)
        		`uvm_info(get_type_name(),$sformatf(" Value of B = %0d", seq.B),UVM_LOW)
            `uvm_info(get_type_name(),$sformatf(" Value of A nor B = %0d", seq.Result),UVM_LOW)
        		$display("-----------------------------------------------------------------------------");
      			end
     	 		else begin
        		`uvm_info(get_type_name(),$sformatf(" TEST FAILED  "),UVM_LOW)
        		end
       			end

       else begin
       //  (seq.Result==8'bX) begin
          `uvm_info(get_type_name(),$sformatf(" DEFAULT VALUE IS INITIATED  "),UVM_LOW)
        end
      
      
        end
  endtask : run_phase
endclass : scoreboard
      
        		